LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE processor_pack IS

CONSTANT NBIT		: INTEGER:=32;
CONSTANT NBYTE	: INTEGER:=8;
CONSTANT NSEL		: INTEGER:=5;

CONSTANT rs_default 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
CONSTANT rt_default 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
CONSTANT rd_default 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
CONSTANT shift_amou		: STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
CONSTANT so_default		: STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');

CONSTANT R_opcode : STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
CONSTANT J_opcode : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000100";
-- CONSTANT L_opcode : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100011";
-- CONSTANT S_opcode : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101011";

END processor_pack;
